* Sample PEX circuit
* Not a complete netlist. Do not use for real simulation.
* This file is only intended for use in testing Substrate's parsers.
* Copyright 2024, Rahul Kumar. All rights reserved.
* 
.subckt sram22_512x64m4w8  VSS VDD ADDR[8] CLK ADDR[7] ADDR[6] ADDR[5] ADDR[4]
+ ADDR[3] ADDR[2] ADDR[1] ADDR[0] WE WMASK[0] DIN[0] DIN[1] DIN[2] DIN[3] DIN[4]
+ DIN[5] DIN[6] DIN[7] WMASK[1] DIN[8] DIN[9] DIN[10] DIN[11] DIN[12] DIN[13]
+ DIN[14] DIN[15] WMASK[2] DIN[16] DIN[17] DIN[18] DIN[19] DIN[20] DIN[21]
+ DIN[22] DIN[23] WMASK[3] DIN[24] DIN[25] DIN[26] DIN[27] DIN[28] DIN[29]
+ DIN[30] DIN[31] WMASK[4] DIN[32] DIN[33] DIN[34] DIN[35] DIN[36] DIN[37]
+ DIN[38] DIN[39] WMASK[5] DIN[40] DIN[41] DIN[42] DIN[43] DIN[44] DIN[45]
+ DIN[46] DIN[47] WMASK[6] DIN[48] DIN[49] DIN[50] DIN[51] DIN[52] DIN[53]
+ DIN[54] DIN[55] WMASK[7] DIN[56] DIN[57] DIN[58] DIN[59] DIN[60] DIN[61]
+ DIN[62] DIN[63] DOUT[0] DOUT[1] DOUT[2] DOUT[3] DOUT[4] DOUT[5] DOUT[6]
+ DOUT[7] DOUT[8] DOUT[9] DOUT[10] DOUT[11] DOUT[12] DOUT[13] DOUT[14] DOUT[15]
+ DOUT[16] DOUT[17] DOUT[18] DOUT[19] DOUT[20] DOUT[21] DOUT[22] DOUT[23]
+ DOUT[24] DOUT[25] DOUT[26] DOUT[27] DOUT[28] DOUT[29] DOUT[30] DOUT[31]
+ DOUT[32] DOUT[33] DOUT[34] DOUT[35] DOUT[36] DOUT[37] DOUT[38] DOUT[39]
+ DOUT[40] DOUT[41] DOUT[42] DOUT[43] DOUT[44] DOUT[45] DOUT[46] DOUT[47]
+ DOUT[48] DOUT[49] DOUT[50] DOUT[51] DOUT[52] DOUT[53] DOUT[54] DOUT[55]
+ DOUT[56] DOUT[57] DOUT[58] DOUT[59] DOUT[60] DOUT[61] DOUT[62] DOUT[63]
* 
* DOUT[63]	DOUT[63]
* DOUT[62]	DOUT[62]
* DOUT[61]	DOUT[61]
* DOUT[60]	DOUT[60]
* DOUT[59]	DOUT[59]
* DOUT[58]	DOUT[58]
* DOUT[57]	DOUT[57]
* DOUT[56]	DOUT[56]
* DOUT[55]	DOUT[55]
* DOUT[54]	DOUT[54]
MX0/Xreplica_bitcell_array/Xcolend_0_0/X0/X0/M0
+ N_X0/RBR_X0/Xreplica_bitcell_array/Xcolend_0_0/X0/X0/M0_s
+ N_VSS_X0/Xreplica_bitcell_array/Xcolend_0_0/X0/X0/M0_g
+ N_X0/RBR_X0/Xreplica_bitcell_array/Xcolend_0_0/X0/X0/M0_s
+ N_VSS_X0/Xreplica_bitcell_array/Xcolend_0_0/X0/X0/M0_b NPASS L=0.14 W=0.14
+ AD=0.0084 AS=0.0084 PD=0.19 PS=0.19 NRD=0 NRS=0 M=1 R=1 SA=0.0602 SB=0.0602
+ UDEF_A=0.0196 UDEF_P=0.56 MULT=1
MX0/Xbitcell_array/Xdummy_col_right_129/X0/X6/M0
+ N_X0/XBITCELL_ARRAY/XDUMMY_COL_RIGHT_129/X0/Q_X0/Xbitcell_array/Xdummy_col_right_129/X0/X3/M0_s
+ N_X0/XBITCELL_ARRAY/XDUMMY_COL_RIGHT_129/X0/QB_X0/Xbitcell_array/Xdummy_col_right_129/X0/X6/M0_g
+ N_VDD_X0/Xbitcell_array/Xdummy_col_right_129/X0/X5/M0_d
+ N_VDD_X0/Xaddr_we_dffs/Xdff_8/X0/X2/M0_b PPU L=0.15 W=0.14 AD=0.0175 AS=0.0428
+ PD=0.39 PS=0.705 NRD=0 NRS=352.788 M=1 R=0.933333 SA=75000.6 SB=75000.2
+ A=0.021 P=0.58 MULT=1
DX285977_noxref noxref_1 N_VDD_X0/Xaddr_we_dffs/Xdff_8/X0/X2/M0_b NWDIODE
+ A=78.8112 P=0
DX285978_noxref noxref_1 N_VDD_X0/Xaddr_we_dffs/Xdff_8/X0/X2/M0_b DNWDIODE_PSUB
+ A=241797 P=1966.92
DX285979_noxref N_VSS_X0/Xreplica_bitcell_array/Xcolend_0_0/X0/X0/M0_b
+ N_VDD_X0/Xaddr_we_dffs/Xdff_8/X0/X2/M0_b DNWDIODE_PW A=188134 P=70753.3
c_1 X0/XADDR_WE_DFFS/XDFF_8/X0/A_197_712# 0 0.0274883f $X=-71.055 $Y=-228.54
c_2 X0/XADDR_WE_DFFS/XDFF_8/X0/A_389_712# 0 0.0145293f $X=-70.095 $Y=-228.54
c_3 X0/XADDR_WE_DFFS/XDFF_8/X0/A_547_712# 0 0.0246353f $X=-69.305 $Y=-228.54
c_599 X0/XCOL_CIRCUITRY/XWMASK_DFFS/XDFF_3/X0/A_197_102# 0 0.0094849f $X=150.665
+ $Y=-117.015
c_600 X0/XCOL_CIRCUITRY/XCOL_GROUP_24/XDFF/X0/A_197_102# 0 0.0094849f $X=150.665
+ $Y=-109.31
c_601 X0/XCOL_CIRCUITRY/XCOL_GROUP_25/XDFF/X0/A_197_102# 0 0.0094849f $X=156.765
+ $Y=-109.31
c_602 X0/XCOL_CIRCUITRY/XCOL_GROUP_26/XDFF/X0/A_197_102# 0 0.0094849f $X=162.865
+ $Y=-109.31
*
.ends
*
*
