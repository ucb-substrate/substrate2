* inverter

.subckt resistor pos neg
R0 pos neg 100
.ends
