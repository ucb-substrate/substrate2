* GENERATED FILE
{% for path in source_paths %}
.include {{path}}
{% endfor %}
