* voltage divider with duplicate subcircuits

.include res_100.spice
.include res_200.spice

.subckt vdivider pwr_vdd pwr_vss out
Rtop pwr_vdd out 600
Xbot out pwr_vss resistor
.ends
