* CMOS buffer

.subckt buffer din dout vdd vss
X0 din dinb vdd vss inverter
X1 dinb dout vdd vss inverter
.ends

.subckt inverter din dout vdd vss
X0 dout din vss vss nshort w=2 l=0.15
X1 dout din vdd vdd pshort w=4 l=0.15
.ends
